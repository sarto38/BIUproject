
`include "AND.v"
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:56:05 01/14/2020 
// Design Name: 
// Module Name:    AND_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module AND_tb();
wire[2:0] out;
reg[2:0] inb, ina;
reg[2:0] rin;
reg clk = 1'b0;
reg AndEnable;
wire AndDone;
AND #(.D(3)) my_gate ( .ina(ina), .inb(inb) ,.rin(rin) ,.AndEnable(AndEnable),.AndDone(AndDone), .out(out), .clk(clk) );

always #1 clk = ~clk;

initial
begin

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b000;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b001;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b010;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b011;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b100;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b101;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b110;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b000;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b001;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b010;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b011;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b100;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b101;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b110;
rin = 3'b111;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b000;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b001;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b010;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b011;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b100;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b101;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b110;

#1
AndEnable= 1'b1;
#6
//////////////////////////////////////////////////////////////////////////////////
    

AndEnable= 1'b0;
#1

ina = 3'b111;
inb = 3'b111;
rin = 3'b111;

#1
AndEnable= 1'b1;


end


endmodule
